module GeradorImm(
    input clock,
    input [12:0] imediato,
    output reg [31:0] imm_estendido,
);

endmodule